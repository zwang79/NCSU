package emu_type_pkg;

typedef enum bit [1:0] {UNKNOWN, READ, WRITE} i2c_op_t;

endpackage
